
module ParallelPrefixCircuit(outputflag, inputflag);

input [65:0] inputflag;
output [65:0] outputflag;
wire [65:0] output1;
wire [65:0] output2;
wire [65:0] output3;
wire [65:0] output4;
wire [65:0] output5;

assign output1[65:64] = (^inputflag[65:64]) ? {inputflag[63],inputflag[62]} : inputflag[65:64];
assign output1[63:62] = (^inputflag[63:62]) ? {inputflag[61],inputflag[60]} : inputflag[63:62];
assign output1[61:60] = (^inputflag[61:60]) ? {inputflag[59],inputflag[58]} : inputflag[61:60];
assign output1[59:58] = (^inputflag[59:58]) ? {inputflag[57],inputflag[56]} : inputflag[59:58];
assign output1[57:56] = (^inputflag[57:56]) ? {inputflag[55],inputflag[54]} : inputflag[57:56];
assign output1[55:54] = (^inputflag[55:54]) ? {inputflag[53],inputflag[52]} : inputflag[55:54];
assign output1[53:52] = (^inputflag[53:52]) ? {inputflag[51],inputflag[50]} : inputflag[53:52];
assign output1[51:50] = (^inputflag[51:50]) ? {inputflag[49],inputflag[48]} : inputflag[51:50];
assign output1[49:48] = (^inputflag[49:48]) ? {inputflag[47],inputflag[46]} : inputflag[49:48];
assign output1[47:46] = (^inputflag[47:46]) ? {inputflag[45],inputflag[44]} : inputflag[47:46];
assign output1[45:44] = (^inputflag[45:44]) ? {inputflag[43],inputflag[42]} : inputflag[45:44];
assign output1[43:42] = (^inputflag[43:42]) ? {inputflag[41],inputflag[40]} : inputflag[43:42];
assign output1[41:40] = (^inputflag[41:40]) ? {inputflag[39],inputflag[38]} : inputflag[41:40];
assign output1[39:38] = (^inputflag[39:38]) ? {inputflag[37],inputflag[36]} : inputflag[39:38];
assign output1[37:36] = (^inputflag[37:36]) ? {inputflag[35],inputflag[34]} : inputflag[37:36];
assign output1[35:34] = (^inputflag[35:34]) ? {inputflag[33],inputflag[32]} : inputflag[35:34];
assign output1[33:32] = (^inputflag[33:32]) ? {inputflag[31],inputflag[30]} : inputflag[33:32];
assign output1[31:30] = (^inputflag[31:30]) ? {inputflag[29],inputflag[28]} : inputflag[31:30];
assign output1[29:28] = (^inputflag[29:28]) ? {inputflag[27],inputflag[26]} : inputflag[29:28];
assign output1[27:26] = (^inputflag[27:26]) ? {inputflag[25],inputflag[24]} : inputflag[27:26];
assign output1[25:24] = (^inputflag[25:24]) ? {inputflag[23],inputflag[22]} : inputflag[25:24];
assign output1[23:22] = (^inputflag[23:22]) ? {inputflag[21],inputflag[20]} : inputflag[23:22];
assign output1[21:20] = (^inputflag[21:20]) ? {inputflag[19],inputflag[18]} : inputflag[21:20];
assign output1[19:18] = (^inputflag[19:18]) ? {inputflag[17],inputflag[16]} : inputflag[19:18];
assign output1[17:16] = (^inputflag[17:16]) ? {inputflag[15],inputflag[14]} : inputflag[17:16];
assign output1[15:14] = (^inputflag[15:14]) ? {inputflag[13],inputflag[12]} : inputflag[15:14];
assign output1[13:12] = (^inputflag[13:12]) ? {inputflag[11],inputflag[10]} : inputflag[13:12];
assign output1[11:10] = (^inputflag[11:10]) ? {inputflag[9],inputflag[8]} : inputflag[11:10];
assign output1[9:8] = (^inputflag[9:8]) ? {inputflag[7],inputflag[6]} : inputflag[9:8];
assign output1[7:6] = (^inputflag[7:6]) ? {inputflag[5],inputflag[4]} : inputflag[7:6];
assign output1[5:4] = (^inputflag[5:4]) ? {inputflag[3],inputflag[2]} : inputflag[5:4];
assign output1[3:2] = (^inputflag[3:2]) ? {inputflag[1],inputflag[0]} : inputflag[3:2];
assign output1[1:0] = inputflag[1:0];

assign output2[65:64] = (^output1[65:64]) ? {output1[61],output1[60]} : output1[65:64];
assign output2[63:62] = (^output1[63:62]) ? {output1[59],output1[58]} : output1[63:62];
assign output2[61:60] = (^output1[61:60]) ? {output1[57],output1[56]} : output1[61:60];
assign output2[59:58] = (^output1[59:58]) ? {output1[55],output1[54]} : output1[59:58];
assign output2[57:56] = (^output1[57:56]) ? {output1[53],output1[52]} : output1[57:56];
assign output2[55:54] = (^output1[55:54]) ? {output1[51],output1[50]} : output1[55:54];
assign output2[53:52] = (^output1[53:52]) ? {output1[49],output1[48]} : output1[53:52];
assign output2[51:50] = (^output1[51:50]) ? {output1[47],output1[46]} : output1[51:50];
assign output2[49:48] = (^output1[49:48]) ? {output1[45],output1[44]} : output1[49:48];
assign output2[47:46] = (^output1[47:46]) ? {output1[43],output1[42]} : output1[47:46];
assign output2[45:44] = (^output1[45:44]) ? {output1[41],output1[40]} : output1[45:44];
assign output2[43:42] = (^output1[43:42]) ? {output1[39],output1[38]} : output1[43:42];
assign output2[41:40] = (^output1[41:40]) ? {output1[37],output1[36]} : output1[41:40];
assign output2[39:38] = (^output1[39:38]) ? {output1[35],output1[34]} : output1[39:38];
assign output2[37:36] = (^output1[37:36]) ? {output1[33],output1[32]} : output1[37:36];
assign output2[35:34] = (^output1[35:34]) ? {output1[31],output1[30]} : output1[35:34];
assign output2[33:32] = (^output1[33:32]) ? {output1[29],output1[28]} : output1[33:32];
assign output2[31:30] = (^output1[31:30]) ? {output1[27],output1[26]} : output1[31:30];
assign output2[29:28] = (^output1[29:28]) ? {output1[25],output1[24]} : output1[29:28];
assign output2[27:26] = (^output1[27:26]) ? {output1[23],output1[22]} : output1[27:26];
assign output2[25:24] = (^output1[25:24]) ? {output1[21],output1[20]} : output1[25:24];
assign output2[23:22] = (^output1[23:22]) ? {output1[19],output1[18]} : output1[23:22];
assign output2[21:20] = (^output1[21:20]) ? {output1[17],output1[16]} : output1[21:20];
assign output2[19:18] = (^output1[19:18]) ? {output1[15],output1[14]} : output1[19:18];
assign output2[17:16] = (^output1[17:16]) ? {output1[13],output1[12]} : output1[17:16];
assign output2[15:14] = (^output1[15:14]) ? {output1[11],output1[10]} : output1[15:14];
assign output2[13:12] = (^output1[13:12]) ? {output1[9],output1[8]} : output1[13:12];
assign output2[11:10] = (^output1[11:10]) ? {output1[7],output1[6]} : output1[11:10];
assign output2[9:8] = (^output1[9:8]) ? {output1[5],output1[4]} : output1[9:8];
assign output2[7:6] = (^output1[7:6]) ? {output1[3],output1[2]} : output1[7:6];
assign output2[5:4] = (^output1[5:4]) ? {output1[1],output1[0]} : output1[5:4];
assign output2[3:0] = output1[3:0];

assign output3[65:64] = (^output2[65:64]) ? {output2[57],output2[56]} : output2[65:64];
assign output3[63:62] = (^output2[63:62]) ? {output2[55],output2[54]} : output2[63:62];
assign output3[61:60] = (^output2[61:60]) ? {output2[53],output2[52]} : output2[61:60];
assign output3[59:58] = (^output2[59:58]) ? {output2[51],output2[50]} : output2[59:58];
assign output3[57:56] = (^output2[57:56]) ? {output2[49],output2[48]} : output2[57:56];
assign output3[55:54] = (^output2[55:54]) ? {output2[47],output2[46]} : output2[55:54];
assign output3[53:52] = (^output2[53:52]) ? {output2[45],output2[44]} : output2[53:52];
assign output3[51:50] = (^output2[51:50]) ? {output2[43],output2[42]} : output2[51:50];
assign output3[49:48] = (^output2[49:48]) ? {output2[41],output2[40]} : output2[49:48];
assign output3[47:46] = (^output2[47:46]) ? {output2[39],output2[38]} : output2[47:46];
assign output3[45:44] = (^output2[45:44]) ? {output2[37],output2[36]} : output2[45:44];
assign output3[43:42] = (^output2[43:42]) ? {output2[35],output2[34]} : output2[43:42];
assign output3[41:40] = (^output2[41:40]) ? {output2[33],output2[32]} : output2[41:40];
assign output3[39:38] = (^output2[39:38]) ? {output2[31],output2[30]} : output2[39:38];
assign output3[37:36] = (^output2[37:36]) ? {output2[29],output2[28]} : output2[37:36];
assign output3[35:34] = (^output2[35:34]) ? {output2[27],output2[26]} : output2[35:34];
assign output3[33:32] = (^output2[33:32]) ? {output2[25],output2[24]} : output2[33:32];
assign output3[31:30] = (^output2[31:30]) ? {output2[23],output2[22]} : output2[31:30];
assign output3[29:28] = (^output2[29:28]) ? {output2[21],output2[20]} : output2[29:28];
assign output3[27:26] = (^output2[27:26]) ? {output2[19],output2[18]} : output2[27:26];
assign output3[25:24] = (^output2[25:24]) ? {output2[17],output2[16]} : output2[25:24];
assign output3[23:22] = (^output2[23:22]) ? {output2[15],output2[14]} : output2[23:22];
assign output3[21:20] = (^output2[21:20]) ? {output2[13],output2[12]} : output2[21:20];
assign output3[19:18] = (^output2[19:18]) ? {output2[11],output2[10]} : output2[19:18];
assign output3[17:16] = (^output2[17:16]) ? {output2[9],output2[8]} : output2[17:16];
assign output3[15:14] = (^output2[15:14]) ? {output2[7],output2[6]} : output2[15:14];
assign output3[13:12] = (^output2[13:12]) ? {output2[5],output2[4]} : output2[13:12];
assign output3[11:10] = (^output2[11:10]) ? {output2[3],output2[2]} : output2[11:10];
assign output3[9:8] = (^output2[9:8]) ? {output2[1],output2[0]} : output2[9:8];
assign output3[7:0] = output2[7:0];

assign output4[65:64] = (^output3[65:64]) ? {output3[49],output3[48]} : output3[65:64];
assign output4[63:62] = (^output3[63:62]) ? {output3[47],output3[46]} : output3[63:62];
assign output4[61:60] = (^output3[61:60]) ? {output3[45],output3[44]} : output3[61:60];
assign output4[59:58] = (^output3[59:58]) ? {output3[43],output3[42]} : output3[59:58];
assign output4[57:56] = (^output3[57:56]) ? {output3[41],output3[40]} : output3[57:56];
assign output4[55:54] = (^output3[55:54]) ? {output3[39],output3[38]} : output3[55:54];
assign output4[53:52] = (^output3[53:52]) ? {output3[37],output3[36]} : output3[53:52];
assign output4[51:50] = (^output3[51:50]) ? {output3[35],output3[34]} : output3[51:50];
assign output4[49:48] = (^output3[49:48]) ? {output3[33],output3[32]} : output3[49:48];
assign output4[47:46] = (^output3[47:46]) ? {output3[31],output3[30]} : output3[47:46];
assign output4[45:44] = (^output3[45:44]) ? {output3[29],output3[28]} : output3[45:44];
assign output4[43:42] = (^output3[43:42]) ? {output3[27],output3[26]} : output3[43:42];
assign output4[41:40] = (^output3[41:40]) ? {output3[25],output3[24]} : output3[41:40];
assign output4[39:38] = (^output3[39:38]) ? {output3[23],output3[22]} : output3[39:38];
assign output4[37:36] = (^output3[37:36]) ? {output3[21],output3[20]} : output3[37:36];
assign output4[35:34] = (^output3[35:34]) ? {output3[19],output3[18]} : output3[35:34];
assign output4[33:32] = (^output3[33:32]) ? {output3[17],output3[16]} : output3[33:32];
assign output4[31:30] = (^output3[31:30]) ? {output3[15],output3[14]} : output3[31:30];
assign output4[29:28] = (^output3[29:28]) ? {output3[13],output3[12]} : output3[29:28];
assign output4[27:26] = (^output3[27:26]) ? {output3[11],output3[10]} : output3[27:26];
assign output4[25:24] = (^output3[25:24]) ? {output3[9],output3[8]} : output3[25:24];
assign output4[23:22] = (^output3[23:22]) ? {output3[7],output3[6]} : output3[23:22];
assign output4[21:20] = (^output3[21:20]) ? {output3[5],output3[4]} : output3[21:20];
assign output4[19:18] = (^output3[19:18]) ? {output3[3],output3[2]} : output3[19:18];
assign output4[17:16] = (^output3[17:16]) ? {output3[1],output3[0]} : output3[17:16];
assign output4[15:0] = output3[15:0];

assign output5[65:64] = (^output4[65:64]) ? {output4[33],output4[32]} : output4[65:64];
assign output5[63:62] = (^output4[63:62]) ? {output4[31],output4[30]} : output4[63:62];
assign output5[61:60] = (^output4[61:60]) ? {output4[29],output4[28]} : output4[61:60];
assign output5[59:58] = (^output4[59:58]) ? {output4[27],output4[26]} : output4[59:58];
assign output5[57:56] = (^output4[57:56]) ? {output4[25],output4[24]} : output4[57:56];
assign output5[55:54] = (^output4[55:54]) ? {output4[23],output4[22]} : output4[55:54];
assign output5[53:52] = (^output4[53:52]) ? {output4[21],output4[20]} : output4[53:52];
assign output5[51:50] = (^output4[51:50]) ? {output4[19],output4[18]} : output4[51:50];
assign output5[49:48] = (^output4[49:48]) ? {output4[17],output4[16]} : output4[49:48];
assign output5[47:46] = (^output4[47:46]) ? {output4[15],output4[14]} : output4[47:46];
assign output5[45:44] = (^output4[45:44]) ? {output4[13],output4[12]} : output4[45:44];
assign output5[43:42] = (^output4[43:42]) ? {output4[11],output4[10]} : output4[43:42];
assign output5[41:40] = (^output4[41:40]) ? {output4[9],output4[8]} : output4[41:40];
assign output5[39:38] = (^output4[39:38]) ? {output4[7],output4[6]} : output4[39:38];
assign output5[37:36] = (^output4[37:36]) ? {output4[5],output4[4]} : output4[37:36];
assign output5[35:34] = (^output4[35:34]) ? {output4[3],output4[2]} : output4[35:34];
assign output5[33:32] = (^output4[33:32]) ? {output4[1],output4[0]} : output4[33:32];
assign output5[31:0] = output4[31:0];

assign outputflag[65:64] = (^output5[65:64]) ? {output5[1],output5[0]} : output5[65:64];
assign outputflag[63:0] = output5[63:0];

endmodule
