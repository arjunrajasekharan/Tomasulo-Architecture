

module CSA1 (a1, a2, a3, b1, b2); // 32 X 33 x 34 -> 34 x 34

input [31:0] a1;
input [32:0] a2;
input [33:0] a3;
output [33:0] b1;
output [33:0] b2;

fullAdder FA1(a1[0], a2[0], a3[0], b1[0], b2[1]);
fullAdder FA2(a1[1], a2[1], a3[1], b1[1], b2[2]);
fullAdder FA3(a1[2], a2[2], a3[2], b1[2], b2[3]);
fullAdder FA4(a1[3], a2[3], a3[3], b1[3], b2[4]);
fullAdder FA5(a1[4], a2[4], a3[4], b1[4], b2[5]);
fullAdder FA6(a1[5], a2[5], a3[5], b1[5], b2[6]);
fullAdder FA7(a1[6], a2[6], a3[6], b1[6], b2[7]);
fullAdder FA8(a1[7], a2[7], a3[7], b1[7], b2[8]);
fullAdder FA9(a1[8], a2[8], a3[8], b1[8], b2[9]);
fullAdder FA10(a1[9], a2[9], a3[9], b1[9], b2[10]);

fullAdder FA11(a1[10], a2[10], a3[10], b1[10], b2[11]);
fullAdder FA12(a1[11], a2[11], a3[11], b1[11], b2[12]);
fullAdder FA13(a1[12], a2[12], a3[12], b1[12], b2[13]);
fullAdder FA14(a1[13], a2[13], a3[13], b1[13], b2[14]);
fullAdder FA15(a1[14], a2[14], a3[14], b1[14], b2[15]);
fullAdder FA16(a1[15], a2[15], a3[15], b1[15], b2[16]);
fullAdder FA17(a1[16], a2[16], a3[16], b1[16], b2[17]);
fullAdder FA18(a1[17], a2[17], a3[17], b1[17], b2[18]);
fullAdder FA19(a1[18], a2[18], a3[18], b1[18], b2[19]);
fullAdder FA20(a1[19], a2[19], a3[19], b1[19], b2[20]);

fullAdder FA21(a1[20], a2[20], a3[20], b1[20], b2[21]);
fullAdder FA22(a1[21], a2[21], a3[21], b1[21], b2[22]);
fullAdder FA23(a1[22], a2[22], a3[22], b1[22], b2[23]);
fullAdder FA24(a1[23], a2[23], a3[23], b1[23], b2[24]);
fullAdder FA25(a1[24], a2[24], a3[24], b1[24], b2[25]);
fullAdder FA26(a1[25], a2[25], a3[25], b1[25], b2[26]);
fullAdder FA27(a1[26], a2[26], a3[26], b1[26], b2[27]);
fullAdder FA28(a1[27], a2[27], a3[27], b1[27], b2[28]);
fullAdder FA29(a1[28], a2[28], a3[28], b1[28], b2[29]);
fullAdder FA30(a1[29], a2[29], a3[29], b1[29], b2[30]);

fullAdder FA31(a1[30], a2[30], a3[30], b1[30], b2[31]);
fullAdder FA32(a1[31], a2[31], a3[31], b1[31], b2[32]);
fullAdder FA33(1'b0, a2[32], a3[32], b1[32], b2[33]);

assign b1[33] = a3[33];
assign b2[0] = 1'b0;

endmodule
