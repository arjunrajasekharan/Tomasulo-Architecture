module PPG(res, a, b);

input [31:0] a;
input b;
output [31:0] res;

and and0(res[0], a[0], b);
and and1(res[1], a[1], b);
and and2(res[2], a[2], b);
and and3(res[3], a[3], b);
and and4(res[4], a[4], b);
and and5(res[5], a[5], b);
and and6(res[6], a[6], b);
and and7(res[7], a[7], b);

and and8(res[8], a[8], b);
and and9(res[9], a[9], b);
and and10(res[10], a[10], b);
and and11(res[11], a[11], b);
and and12(res[12], a[12], b);
and and13(res[13], a[13], b);
and and14(res[14], a[14], b);
and and15(res[15], a[15], b);

and and16(res[16], a[16], b);
and and17(res[17], a[17], b);
and and18(res[18], a[18], b);
and and19(res[19], a[19], b);
and and20(res[20], a[20], b);
and and21(res[21], a[21], b);
and and22(res[22], a[22], b);
and and23(res[23], a[23], b);

and and24(res[24], a[24], b);
and and25(res[25], a[25], b);
and and26(res[26], a[26], b);
and and27(res[27], a[27], b);
and and28(res[28], a[28], b);
and and29(res[29], a[29], b);
and and30(res[30], a[30], b);
and and31(res[31], a[31], b);

endmodule
